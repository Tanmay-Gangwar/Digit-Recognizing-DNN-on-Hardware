library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all;

entity dataType_tb is
end entity;

architecture Behavioral of dataType_tb is
    begin
    end Behavioral;